* Extracted by KLayout with SG13G2 LVS runset on : 30/04/2024 14:49

* cell rdiv_notsep
.SUBCKT rdiv_notsep
* device instance $1 r0 *1 2.272,-22.301 res_rhigh
R$1 IN_P \$3 res_rhigh w=0.5 l=15.0 b=0.0 ps=0.0 m=1.0
* device instance $2 r0 *1 4.292,-14.879 res_rhigh
R$2 \$2 \$3 res_rhigh w=0.5 l=7.5 b=0.0 ps=0.0 m=1.0
* device instance $3 r0 *1 6.681,-14.879 res_rhigh
R$3 \$2 \$4 res_rhigh w=0.5 l=7.5 b=0.0 ps=0.0 m=1.0
* device instance $4 r0 *1 -0.987,-10.023 res_rhigh
R$4 IN_P VOUT res_rhigh w=0.5 l=10.0 b=0.0 ps=0.0 m=1.0
.ENDS rdiv_notsep
