* Extracted by KLayout with SG13G2 LVS runset on : 30/04/2024 10:13

* cell nmos_current_mirror
* pin VS
* pin VOUT
* pin IREF
* pin VSS
.SUBCKT nmos_current_mirror VS VOUT IREF VSS
* device instance $1 r0 *1 0.736,1.102 sg13_lv_nmos
M$1 VS IREF VSS VSS sg13_lv_nmos W=6.0 L=2.0
* device instance $2 r0 *1 3.116,1.102 sg13_lv_nmos
M$2 VSS IREF VOUT VSS sg13_lv_nmos W=24.0 L=2.0
* device instance $6 r0 *1 12.636,1.102 sg13_lv_nmos
M$6 VSS IREF IREF VSS sg13_lv_nmos W=6.0 L=2.0
.ENDS nmos_current_mirror
