* Extracted by KLayout with SG13G2 LVS runset on : 30/04/2024 10:34

* cell OTA_without_rcomp
* pin VOUT
* pin VMID2
* pin VSS
* pin VS
* pin IREF
* pin VDD
* pin VMID1
* pin VIN_P
* pin VIN_N
* pin sub!
.SUBCKT OTA_without_rcomp VOUT VMID2 VSS VS IREF VDD VMID1 VIN_P VIN_N sub!
* device instance $1 r0 *1 -28.27,-7.193 sg13_lv_nmos
M$1 VS IREF VSS sub! sg13_lv_nmos W=6.0 L=2.0
* device instance $2 r0 *1 -25.89,-7.193 sg13_lv_nmos
M$2 VSS IREF VOUT sub! sg13_lv_nmos W=24.0 L=2.0
* device instance $6 r0 *1 -16.37,-7.193 sg13_lv_nmos
M$6 VSS IREF IREF sub! sg13_lv_nmos W=6.0 L=2.0
* device instance $13 r0 *1 -10.772,3.507 sg13_lv_nmos
M$13 VMID1 VIN_N VS sub! sg13_lv_nmos W=15.0 L=2.0
* device instance $14 r0 *1 -8.392,3.507 sg13_lv_nmos
M$14 VS VIN_P VMID2 sub! sg13_lv_nmos W=15.0 L=2.0
* device instance $21 r0 *1 8.788,-1.299 sg13_lv_pmos
M$21 VDD VMID2 VOUT \$19 sg13_lv_pmos W=20.0 L=0.5
* device instance $29 r0 *1 -9.278,14.481 sg13_lv_pmos
M$29 VMID2 VMID1 VDD \$19 sg13_lv_pmos W=2.0 L=1.0
* device instance $30 r0 *1 -7.898,14.481 sg13_lv_pmos
M$30 VDD VMID1 VMID1 \$19 sg13_lv_pmos W=2.0 L=1.0
* device instance $33 r0 *1 -26.07,-57.903 cap_cmim
C$33 VOUT VMID2 cap_cmim w=45 l=45 m=1
.ENDS OTA_without_rcomp
