* Extracted by KLayout with SG13G2 LVS runset on : 29/04/2024 13:56

* cell TOP
.SUBCKT TOP
* device instance $1 r0 *1 14.014,3.8 res_rhigh
R$1 \$1 \$2 res_rhigh w=0.5 l=2.5 b=0.0 ps=0.0 m=1.0
* device instance $2 r0 *1 17.047,8.495 res_rhigh
R$2 \$2 \$3 res_rhigh w=0.5 l=2.5 b=0.0 ps=0.0 m=1.0
* device instance $3 r0 *1 15.525,13.191 res_rhigh
R$3 \$3 \$4 res_rhigh w=0.5 l=2.5 b=0.0 ps=0.0 m=1.0
* device instance $4 r0 *1 18.544,17.895 res_rhigh
R$4 \$4 \$5 res_rhigh w=0.5 l=2.5 b=0.0 ps=0.0 m=1.0
.ENDS TOP
