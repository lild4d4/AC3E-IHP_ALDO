* Extracted by KLayout with SG13G2 LVS runset on : 30/04/2024 10:21

* cell nmos_diffpar
* pin VS
* pin VMID2
* pin VMID1
* pin VIN_P
* pin VIN_N
* pin VSS
.SUBCKT nmos_diffpar VS VMID2 VMID1 VIN_P VIN_N VSS
* device instance $1 r0 *1 0.865,-3.18 sg13_lv_nmos
M$1 VMID1 VIN_N VS VSS sg13_lv_nmos W=15.0 L=2.0
* device instance $2 r0 *1 3.245,-3.18 sg13_lv_nmos
M$2 VS VIN_P VMID2 VSS sg13_lv_nmos W=15.0 L=2.0
.ENDS nmos_diffpar
