* Extracted by KLayout with SG13G2 LVS runset on : 29/04/2024 17:12

* cell rdiv
* pin IN_P
.SUBCKT rdiv IN_P
* device instance $1 r0 *1 14.024,3.799 res_rhigh
R$1 IN_P \$4 res_rhigh w=0.5 l=5.0 b=0.0 ps=0.0 m=1.0
* device instance $2 r0 *1 15.524,3.799 res_rhigh
R$2 IN_P \$5 res_rhigh w=0.5 l=2.5 b=0.0 ps=0.0 m=1.0
* device instance $4 r0 *1 18.524,3.799 res_rhigh
R$4 \$3 \$2 res_rhigh w=0.5 l=5.0 b=0.0 ps=0.0 m=1.0
* device instance $6 r0 *1 15.524,8.499 res_rhigh
R$6 \$18 \$32 res_rhigh w=0.5 l=5.0 b=0.0 ps=0.0 m=1.0
* device instance $8 r0 *1 18.524,8.499 res_rhigh
R$8 \$3 \$32 res_rhigh w=0.5 l=2.5 b=0.0 ps=0.0 m=1.0
* device instance $9 r0 *1 14.024,13.199 res_rhigh
R$9 \$31 \$47 res_rhigh w=0.5 l=2.5 b=0.0 ps=0.0 m=1.0
* device instance $10 r0 *1 15.524,13.199 res_rhigh
R$10 \$33 \$48 res_rhigh w=0.5 l=5.0 b=0.0 ps=0.0 m=1.0
* device instance $12 r0 *1 18.524,13.199 res_rhigh
R$12 \$34 \$49 res_rhigh w=0.5 l=5.0 b=0.0 ps=0.0 m=1.0
* device instance $14 r0 *1 15.524,17.899 res_rhigh
R$14 \$50 \$52 res_rhigh w=0.5 l=5.0 b=0.0 ps=0.0 m=1.0
* device instance $15 r0 *1 17.024,17.899 res_rhigh
R$15 \$49 \$52 res_rhigh w=0.5 l=2.5 b=0.0 ps=0.0 m=1.0
.ENDS rdiv
