* Extracted by KLayout with SG13G2 LVS runset on : 30/04/2024 15:06

* cell rdiv_testcase
* pin IN_P
* pin VOUT
.SUBCKT rdiv_testcase IN_P VOUT
* device instance $1 r0 *1 2.272,-22.301 res_rhigh
R$1 IN_P \$4 res_rhigh w=0.5 l=15.0 b=0.0 ps=0.0 m=1.0
* device instance $2 r0 *1 6.681,-15.121 res_rhigh
R$2 \$2 \$3 res_rhigh w=0.5 l=15.0 b=0.0 ps=0.0 m=1.0
* device instance $4 r0 *1 -0.987,-10.023 res_rhigh
R$4 IN_P VOUT res_rhigh w=0.5 l=10.0 b=0.0 ps=0.0 m=1.0
.ENDS rdiv_testcase
