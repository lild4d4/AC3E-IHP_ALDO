* Extracted by KLayout with SG13G2 LVS runset on : 26/04/2024 09:04

* cell rcomp
.SUBCKT rcomp
.ENDS rcomp
